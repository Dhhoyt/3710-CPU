module GPUController(
	input wire [15:0] read_data,
	output wire [15:0] read_address
);

endmodule